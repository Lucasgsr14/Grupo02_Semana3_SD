library verilog;
use verilog.vl_types.all;
entity DEMUX_SUM_vlg_vec_tst is
end DEMUX_SUM_vlg_vec_tst;

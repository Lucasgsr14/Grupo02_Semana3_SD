library verilog;
use verilog.vl_types.all;
entity DEMUX_REG_vlg_vec_tst is
end DEMUX_REG_vlg_vec_tst;
